module alu
#(
  parameter WIDTH=8
 )
 (
  input  wire [      2:0] opcode    ,
  input  wire [WIDTH-1:0] in_a      ,
  input  wire [WIDTH-1:0] in_b      ,
  output wire             a_is_zero ,
  output reg  [WIDTH-1:0] alu_out    
 );
	localparam PASS0=0, PASS1=1, ADD=2, AND=3, XOR=4, PASSB=5, PASS6=6, PASS7=7;
always @*
    case(opcode)
      PASS0, PASS1, PASS6, PASS7: alu_out = in_a;
			ADD  : alu_out = in_a + in_b;
			AND  : alu_out = in_a & in_b;
			XOR  : alu_out = in_a ^ in_b;
			PASSB: alu_out = in_b;
    endcase
assign a_is_zero = (in_a == 0) ? 8'b1 : 0;	
endmodule
